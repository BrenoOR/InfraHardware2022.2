module signext32_16 (
    input wire [15:0] data_input;
    output wire [31:0] data_out;
);

endmodule